module not32bit(out, A);

input [31:0] A; 
output [31:0] out; 

not g0(out[0], A[0] );
not g1(out[1], A[1]); 
not g2(out[2], A[2]);
not g3(out[3], A[3]);
not g4(out[4], A[4]);
not g5(out[5], A[5]);
not g6(out[6], A[6]);
not g7(out[7], A[7]);
not g8(out[8], A[8]);
not g9(out[9], A[9]);
not g10(out[10], A[10]);
not g11(out[11], A[11]);
not g12(out[12], A[12]);
not g13(out[13], A[13]);
not g14(out[14], A[14]);
not g15(out[15], A[15]);
not g16(out[16], A[16]);
not g17(out[17], A[17]);
not g18(out[18], A[18]);
not g19(out[19], A[19]);
not g20(out[20], A[20]);
not g21(out[21], A[21]); 
not g22(out[22], A[22]);
not g23(out[23], A[23]);
not g24(out[24], A[24]);
not g25(out[25], A[25]);
not g26(out[26], A[26]);
not g27(out[27], A[27]);
not g28(out[28], A[28]);
not g29(out[29], A[29]);
not g30(out[30], A[30]);
not g31(out[31], A[31]); 

endmodule 